module part2(SW, KEY, LEDR, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5);
      
		input [9:0] SW;
		input [3:0] KEY;
		input [6:0] HEX0;
		input [6:0] HEX1;
		input [6:0] HEX2;
		input [6:0] HEX3;
		input [6:0] HEX4;
		input [6:0] HEX5;
		output [7:0] LEDR;
		
		wire [7:0] W2;
	   wire [7:0] W3;
		wire [3:0] W4;
		assign W4 = 4'b0000;
		
	   Display U1(.in(SW[3:0]), .out(HEX0[6:0]));
	   ALU U2(.I1(SW[3:0]), .I2(W3[7:0]), .Key(KEY[3:1]), .Out(W2[7:0]));
		Register U3(.Clock(KEY[0]), .Reset_b(SW[9]), .I(W2[7:0]), .O(W3[7:0]));
		
		assign LEDR = W3;
		Display U4(.in(W3[7:4]), .out(HEX4[6:0]));//MSB
		Display U5(.in(W3[3:0]), .out(HEX5[6:0]));//LSB
		Display U6(.in(W4[3:0]), .out(HEX1[6:0]));
		Display U7(.in(W4[3:0]), .out(HEX2[6:0]));
		Display U8(.in(W4[3:0]), .out(HEX3[6:0]));
		
endmodule
 
 
module Register(Clock, Reset_b, I, O);

	  input Clock;
	  input Reset_b;
	  input [7:0] I;
	  output reg [7:0] O; //output
	  always@(posedge Clock)
	  begin
		 if(Reset_b == 1'b0)
		  begin
			O <= 0;
		  end
		 else
		  begin	
			O <= I;
	     end  
	  end
	  
endmodule


module ALU(I1, I2, Key, Out);

     input [7:0] I2;
	  input [3:0] I1;
	  input [3:1] Key;
	  
	  output [7:0] Out;
	 
	  wire[3:0] A, B;
	  wire[7:0] C;
	  assign A = I1 [3:0];
	  assign B = I2 [7:4];
	  assign C = I2 [7:0];
		
	  reg [7:0] ALUout;
	  wire[3:0] w1; //Selector  
	  wire w2;
	  
	  Adder X1(.A(I1[3:0]), .B(I2[7:4]), .Cout(w2), .S(w1[3:0]), .Cin(0));
	  
	  always@(*)
		begin
		  case(Key[3:1])
				
				3'b000: ALUout = {3'b000,w2, w1};
				
				3'b001: ALUout = {4'b0000,A + B};
				
				3'b010: ALUout = {~(A|B),~(A&B)};
				
				3'b011: begin
							 if((|A)||(|B) == 1) //bitwise OR
								ALUout = 8'b11000000;
							 else ALUout = 8'b00000000; 
						  end
				
				3'b100: begin
							 if((A == 4'b0011||4'b0110||4'b1100||4'b1010||4'b0101||4'b1001) && (B == 4'b0111||4'b1110||4'b1011||4'b1101))
								ALUout = 8'b00111111;
							 else ALUout = 8'b00000000;
						  end
				3'b101: 
						  ALUout = {B, ~A};
						  
				3'b110: ALUout = {A^B,A~^B};
				3'b111: ALUout = C;
				default: ALUout = 8'b00000000;
		  endcase
		end
		assign Out = ALUout;
		
endmodule
  
  
module Adder(Cin, A, B, S, Cout);
  
	  input [3:0] A, B;
	  input Cin;
	  output [3:0] S;
	  output Cout;
	  wire [2:0] W;
	  
	  FullAdd x1(.cin(Cin), .a(A[3]), .b(B[3]), .cout(W[0]), .s(S[3]));    //bit0
	  FullAdd x2(.cin(W[0]), .a(A[2]), .b(B[2]), .cout(W[1]), .s(S[2]));   //bit1
	  FullAdd x3(.cin(W[1]), .a(A[1]), .b(B[1]), .cout(W[2]), .s(S[1]));   //bit2
	  FullAdd x4(.cin(W[2]), .a(A[0]), .b(B[0]), .cout(Cout), .s(S[0]));   //bit3

endmodule

  
module FullAdd(cin, a, b, s, cout);

	  input cin, a, b;
	  output s, cout;
	  assign s = a^b^cin;
	  assign cout = (a&b)|(a&cin)|(b&cin);
	  
endmodule


module Display(in, out); //HEX
  
	 input [3:0] in;
	 reg [6:0] out_wire;
	 output [6:0] out = ~out_wire;
	  
	 always@(*)
	 begin
	 case (in)
		0: out_wire = 7'b0111111;
		1: out_wire = 7'b0000110;
		2: out_wire = 7'b1011011;
		3: out_wire = 7'b1001111;
		4: out_wire = 7'b1100110;
		5: out_wire = 7'b1101101;
		6: out_wire = 7'b1111101;
		7: out_wire = 7'b0000111;
		8: out_wire = 7'b1111111;
		9: out_wire = 7'b1100111;
		10: out_wire = 7'b1110111;
		11: out_wire = 7'b1111100;
		12: out_wire = 7'b0111001;
		13: out_wire = 7'b1011110;
		14: out_wire = 7'b1111001;
		15: out_wire = 7'b1110001;
	 endcase
	 end
	 
endmodule
